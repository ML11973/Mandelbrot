/run/media/leemarc/Shared/Switchdrive/Private/Documents/Master/2_S2/LPSC/Mandelbrot/lpsc-mandelbrot/designs/vivado/lpsc_mandelbrot_firmware/2021.2/src/hdl/lpsc_mandelbrot_firmware.vhd